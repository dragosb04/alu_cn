`ifndef REG_Q_SUB_V
`define REG_Q_SUB_V

module reg_q_sub (
  input CLK, RESET, c1, c2, c4, c6, 
  input [31:0] ibus,
  input a_lsb,
  input sign,
  output reg q_lsb,
  output reg [31:0] obus
);

reg [31:0] q;

always @(posedge CLK, negedge RESET) begin
  if(!RESET)
    q <= 0;
  else if (c1) begin
    q <= ibus;
    q[0] <= 0;
  end else if (c2)
    q[0] <= ~sign;
  else if(c4) 
    begin
        q_lsb <= q[0];
        q <= {q[31], q[31:1]};
        q[31] <= a_lsb;
        q[0] <= 0;
      end

end


always @ (*) begin
  if(c6) 
    obus <= q;
  else obus <= 32'bz;
  
end

endmodule

`endif